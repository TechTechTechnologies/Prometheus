library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity FEEDBACK_CONTROLLER is
  port
  (
    
  );
begin



end;